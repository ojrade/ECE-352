module bin2bcd(
  input 	[3:0] bin,		// can be from 0 to 15
  output	[3:0] upper,	// upper digit as BCD
  output	[3:0] lower		// lower digit as BCD
);

  /////////////////////////////////////////
  // Define any needed internal signals //
  ///////////////////////////////////////
  
  
  ////////////////////////////////////////////////
  // Implement bin2bcd producing lower & upper //
  // with a few verilog data flow statements  //
  /////////////////////////////////////////////
  
  
endmodule
  
  