module msg_ROM(
  input [7:0] addr,			// address of msg character to look up
  output reg [7:0] tx_data	// data to be transmitted
);
  
	/////////////////////////////////////////////
	// big comb block that determines message //
    // byte based on {msg,msg_byte_cnt}      //
	// Generated from a perl script.  Yes   //
	// old people use perl not python.     //
	////////////////////////////////////////  
  	always_comb
	  case (addr)
		8'h0 : tx_data = 8'h45;
		8'h1 : tx_data = 8'h43;
		8'h2 : tx_data = 8'h45;
		8'h3 : tx_data = 8'h33;
		8'h4 : tx_data = 8'h35;
		8'h5 : tx_data = 8'h32;
		8'h6 : tx_data = 8'h20;
		8'h7 : tx_data = 8'h69;
		8'h8 : tx_data = 8'h73;
		8'h9 : tx_data = 8'h20;
		8'ha : tx_data = 8'h67;
		8'hb : tx_data = 8'h72;
		8'hc : tx_data = 8'h65;
		8'hd : tx_data = 8'h61;
		8'he : tx_data = 8'h74;
		8'hf : tx_data = 8'h21;
		8'h10 : tx_data = 8'h45;
		8'h11 : tx_data = 8'h43;
		8'h12 : tx_data = 8'h45;
		8'h13 : tx_data = 8'h33;
		8'h14 : tx_data = 8'h35;
		8'h15 : tx_data = 8'h32;
		8'h16 : tx_data = 8'h20;
		8'h17 : tx_data = 8'h73;
		8'h18 : tx_data = 8'h75;
		8'h19 : tx_data = 8'h63;
		8'h1a : tx_data = 8'h6b;
		8'h1b : tx_data = 8'h73;
		8'h1c : tx_data = 8'h45;
		8'h1d : tx_data = 8'h67;
		8'h1e : tx_data = 8'h67;
		8'h1f : tx_data = 8'h73;
		8'h20 : tx_data = 8'h20;
		8'h21 : tx_data = 8'h47;
		8'h22 : tx_data = 8'h6f;
		8'h23 : tx_data = 8'h21;
		8'h24 : tx_data = 8'h20;
		8'h25 : tx_data = 8'h42;
		8'h26 : tx_data = 8'h75;
		8'h27 : tx_data = 8'h63;
		8'h28 : tx_data = 8'h6b;
		8'h29 : tx_data = 8'h79;
		8'h2a : tx_data = 8'h20;
		8'h2b : tx_data = 8'h47;
		8'h2c : tx_data = 8'h6f;
		8'h2d : tx_data = 8'h21;
		8'h2e : tx_data = 8'h21;
		8'h2f : tx_data = 8'h20;
		8'h30 : tx_data = 8'h54;
		8'h31 : tx_data = 8'h68;
		8'h32 : tx_data = 8'h65;
		8'h33 : tx_data = 8'h51;
		8'h34 : tx_data = 8'h75;
		8'h35 : tx_data = 8'h69;
		8'h36 : tx_data = 8'h63;
		8'h37 : tx_data = 8'h6b;
		8'h38 : tx_data = 8'h42;
		8'h39 : tx_data = 8'h72;
		8'h3a : tx_data = 8'h6f;
		8'h3b : tx_data = 8'h77;
		8'h3c : tx_data = 8'h6e;
		8'h3d : tx_data = 8'h46;
		8'h3e : tx_data = 8'h6f;
		8'h3f : tx_data = 8'h78;
		8'h40 : tx_data = 8'h4a;
		8'h41 : tx_data = 8'h75;
		8'h42 : tx_data = 8'h6d;
		8'h43 : tx_data = 8'h70;
		8'h44 : tx_data = 8'h65;
		8'h45 : tx_data = 8'h64;
		8'h46 : tx_data = 8'h20;
		8'h47 : tx_data = 8'h4f;
		8'h48 : tx_data = 8'h76;
		8'h49 : tx_data = 8'h65;
		8'h4a : tx_data = 8'h72;
		8'h4b : tx_data = 8'h20;
		8'h4c : tx_data = 8'h54;
		8'h4d : tx_data = 8'h68;
		8'h4e : tx_data = 8'h65;
		8'h4f : tx_data = 8'h20;
		8'h50 : tx_data = 8'h4c;
		8'h51 : tx_data = 8'h61;
		8'h52 : tx_data = 8'h7a;
		8'h53 : tx_data = 8'h79;
		8'h54 : tx_data = 8'h20;
		8'h55 : tx_data = 8'h44;
		8'h56 : tx_data = 8'h6f;
		8'h57 : tx_data = 8'h67;
		8'h58 : tx_data = 8'h73;
		8'h59 : tx_data = 8'h20;
		8'h5a : tx_data = 8'h49;
		8'h5b : tx_data = 8'h6e;
		8'h5c : tx_data = 8'h64;
		8'h5d : tx_data = 8'h65;
		8'h5e : tx_data = 8'h65;
		8'h5f : tx_data = 8'h64;
		8'h60 : tx_data = 8'h57;
		8'h61 : tx_data = 8'h68;
		8'h62 : tx_data = 8'h79;
		8'h63 : tx_data = 8'h20;
		8'h64 : tx_data = 8'h64;
		8'h65 : tx_data = 8'h69;
		8'h66 : tx_data = 8'h64;
		8'h67 : tx_data = 8'h20;
		8'h68 : tx_data = 8'h49;
		8'h69 : tx_data = 8'h20;
		8'h6a : tx_data = 8'h61;
		8'h6b : tx_data = 8'h6c;
		8'h6c : tx_data = 8'h6c;
		8'h6d : tx_data = 8'h6f;
		8'h6e : tx_data = 8'h77;
		8'h6f : tx_data = 8'h20;
		8'h70 : tx_data = 8'h66;
		8'h71 : tx_data = 8'h6f;
		8'h72 : tx_data = 8'h72;
		8'h73 : tx_data = 8'h20;
		8'h74 : tx_data = 8'h73;
		8'h75 : tx_data = 8'h6f;
		8'h76 : tx_data = 8'h20;
		8'h77 : tx_data = 8'h6d;
		8'h78 : tx_data = 8'h61;
		8'h79 : tx_data = 8'h6e;
		8'h7a : tx_data = 8'h79;
		8'h7b : tx_data = 8'h20;
		8'h7c : tx_data = 8'h70;
		8'h7d : tx_data = 8'h6f;
		8'h7e : tx_data = 8'h73;
		8'h7f : tx_data = 8'h73;
		8'h80 : tx_data = 8'h69;
		8'h81 : tx_data = 8'h62;
		8'h82 : tx_data = 8'h6c;
		8'h83 : tx_data = 8'h65;
		8'h84 : tx_data = 8'h20;
		8'h85 : tx_data = 8'h6d;
		8'h86 : tx_data = 8'h65;
		8'h87 : tx_data = 8'h73;
		8'h88 : tx_data = 8'h73;
		8'h89 : tx_data = 8'h61;
		8'h8a : tx_data = 8'h67;
		8'h8b : tx_data = 8'h65;
		8'h8c : tx_data = 8'h73;
		8'h8d : tx_data = 8'h3f;
		8'h8e : tx_data = 8'h3f;
		8'h8f : tx_data = 8'h20;
		8'h90 : tx_data = 8'h4e;
		8'h91 : tx_data = 8'h6f;
		8'h92 : tx_data = 8'h77;
		8'h93 : tx_data = 8'h20;
		8'h94 : tx_data = 8'h69;
		8'h95 : tx_data = 8'h73;
		8'h96 : tx_data = 8'h20;
		8'h97 : tx_data = 8'h74;
		8'h98 : tx_data = 8'h68;
		8'h99 : tx_data = 8'h65;
		8'h9a : tx_data = 8'h20;
		8'h9b : tx_data = 8'h74;
		8'h9c : tx_data = 8'h69;
		8'h9d : tx_data = 8'h6d;
		8'h9e : tx_data = 8'h65;
		8'h9f : tx_data = 8'h20;
		8'ha0 : tx_data = 8'h66;
		8'ha1 : tx_data = 8'h6f;
		8'ha2 : tx_data = 8'h72;
		8'ha3 : tx_data = 8'h20;
		8'ha4 : tx_data = 8'h61;
		8'ha5 : tx_data = 8'h6c;
		8'ha6 : tx_data = 8'h6c;
		8'ha7 : tx_data = 8'h20;
		8'ha8 : tx_data = 8'h67;
		8'ha9 : tx_data = 8'h6f;
		8'haa : tx_data = 8'h6f;
		8'hab : tx_data = 8'h64;
		8'hac : tx_data = 8'h20;
		8'had : tx_data = 8'h6d;
		8'hae : tx_data = 8'h65;
		8'haf : tx_data = 8'h6e;
		8'hb0 : tx_data = 8'h74;
		8'hb1 : tx_data = 8'h6f;
		8'hb2 : tx_data = 8'h20;
		8'hb3 : tx_data = 8'h63;
		8'hb4 : tx_data = 8'h6f;
		8'hb5 : tx_data = 8'h6d;
		8'hb6 : tx_data = 8'h65;
		8'hb7 : tx_data = 8'h20;
		8'hb8 : tx_data = 8'h74;
		8'hb9 : tx_data = 8'h6f;
		8'hba : tx_data = 8'h20;
		8'hbb : tx_data = 8'h74;
		8'hbc : tx_data = 8'h68;
		8'hbd : tx_data = 8'h65;
		8'hbe : tx_data = 8'h20;
		8'hbf : tx_data = 8'h20;
		8'hc0 : tx_data = 8'h61;
		8'hc1 : tx_data = 8'h69;
		8'hc2 : tx_data = 8'h64;
		8'hc3 : tx_data = 8'h20;
		8'hc4 : tx_data = 8'h6f;
		8'hc5 : tx_data = 8'h66;
		8'hc6 : tx_data = 8'h20;
		8'hc7 : tx_data = 8'h74;
		8'hc8 : tx_data = 8'h68;
		8'hc9 : tx_data = 8'h65;
		8'hca : tx_data = 8'h69;
		8'hcb : tx_data = 8'h72;
		8'hcc : tx_data = 8'h20;
		8'hcd : tx_data = 8'h20;
		8'hce : tx_data = 8'h20;
		8'hcf : tx_data = 8'h20;
		8'hd0 : tx_data = 8'h63;
		8'hd1 : tx_data = 8'h6f;
		8'hd2 : tx_data = 8'h75;
		8'hd3 : tx_data = 8'h6e;
		8'hd4 : tx_data = 8'h74;
		8'hd5 : tx_data = 8'h72;
		8'hd6 : tx_data = 8'h79;
		8'hd7 : tx_data = 8'h2e;
		8'hd8 : tx_data = 8'h20;
		8'hd9 : tx_data = 8'h20;
		8'hda : tx_data = 8'h20;
		8'hdb : tx_data = 8'h20;
		8'hdc : tx_data = 8'h20;
		8'hdd : tx_data = 8'h20;
		8'hde : tx_data = 8'h20;
		8'hdf : tx_data = 8'h20;
		8'he0 : tx_data = 8'h57;
		8'he1 : tx_data = 8'h68;
		8'he2 : tx_data = 8'h79;
		8'he3 : tx_data = 8'h41;
		8'he4 : tx_data = 8'h72;
		8'he5 : tx_data = 8'h65;
		8'he6 : tx_data = 8'h59;
		8'he7 : tx_data = 8'h6f;
		8'he8 : tx_data = 8'h75;
		8'he9 : tx_data = 8'h53;
		8'hea : tx_data = 8'h74;
		8'heb : tx_data = 8'h69;
		8'hec : tx_data = 8'h6c;
		8'hed : tx_data = 8'h6c;
		8'hee : tx_data = 8'h20;
		8'hef : tx_data = 8'h20;
		8'hf0 : tx_data = 8'h20;
		8'hf1 : tx_data = 8'h54;
		8'hf2 : tx_data = 8'h65;
		8'hf3 : tx_data = 8'h73;
		8'hf4 : tx_data = 8'h74;
		8'hf5 : tx_data = 8'h69;
		8'hf6 : tx_data = 8'h6e;
		8'hf7 : tx_data = 8'h67;
		8'hf8 : tx_data = 8'h20;
		8'hf9 : tx_data = 8'h74;
		8'hfa : tx_data = 8'h68;
		8'hfb : tx_data = 8'h69;
		8'hfc : tx_data = 8'h73;
		8'hfd : tx_data = 8'h3f;
		8'hfe : tx_data = 8'h20;
		8'hff : tx_data = 8'h20;
	  endcase
	  
endmodule